--------------------------------------------------
--	Author:      Renato Noskoski Kissel
--	Created:     Nov 14, 2025
--
--	Project:     Atividade Prática 3 - ULA
--	Description: A<B, saida = 1 se A<B, caso contrário, saida = 0.
--               Este arquivo irá ser usado apenas na divisão, apesar da ULA implementar
--               esta operação, ficaria inviável usar a outra lógica já escrita.
--------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- saida = 1, se A for menor do que B,
-- caso o contrário, saida = 0

entity count_less_than_B is
  generic (
    N : positive := 32 -- número de bits das entradas
  );
  port (
    input_a : in STD_LOGIC_VECTOR(N - 1 downto 0); -- entrada A com N bits com sinal
    input_b : in STD_LOGIC_VECTOR(N - 1 downto 0); -- entrada B com N bits com sinal
    result  : out std_logic -- saída
  );
end count_less_than_B;

architecture behavior of count_less_than_B is
  signal result_subtraction : std_logic_vector(N - 1 downto 0);
  signal overflow           : std_logic;

begin
  subtractor : entity work.subtractor(behavior)
    generic map(N => N)
    port map
    (
      input_a   => std_logic_vector(input_a),
      input_b   => std_logic_vector(input_b),
      result    => result_subtraction,
      carry_out => open,
      overflow  => overflow
    );

  result <= overflow xor result_subtraction(N - 1);
end architecture behavior;